module FPGAPOSMachine(input i,
							output o);

endmodule
